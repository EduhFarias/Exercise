LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL

entity test is
  port(
    clk : in std_logic;
  
  
    o : out std_logic_vector : (7 downto 0)
  );
end test;  

architecture arch of test is
  -- uso de signal ou constant
  begin
  
  --uso de when else, ou uso de with ... select /n ... <= with "..."
  
end arch;
  
  
